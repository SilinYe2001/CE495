`ifndef __GLOBALS__
`define __GLOBALS__
// UVM Globals
localparam int CLOCK_PERIOD = 10;


localparam string RAD_IN_NAME="rad.txt";
localparam string COS_OUT_NAME = "cos.txt";
localparam string SIN_OUT_NAME = "sin.txt";
localparam string COS_CMP_NAME = "cos_cmp.txt";
localparam string SIN_CMP_NAME = "sin_cmp.txt";

`endif
